package DRAM;

import FIFO::*;
import FIFOF::*;
import GetPut::*;
import BRAM::*;
import Vector::*;
import TriState::*;
import RegFile::*;
import FuseTestTypes::*;
import List::*;

(* always_ready, always_enabled *)
interface DRAM_ifc;
    // test
    method Action init_test(MemoryInitT minit);

    // system control
    method Action cs(Bit#(1) cs);
    method Action n_oe(Bit#(1) n_oe);
    method Action n_ce(Bit#(1) n_ce);

    // address bus
    method Action addr(Bit#(14) addr);

    // data bus - output only but still needs to be tristate
    interface Inout#(Bit#(8)) data;
endinterface

//(* synthesize *)
module mkDRAM(DRAM_ifc);
    Wire#(Bit#(1)) cs_in <- mkBypassWire;
    Wire#(Bit#(1)) n_oe_in <- mkBypassWire;
    Wire#(Bit#(1)) n_ce_in <- mkBypassWire;

    RegFile#(Bit#(14), Bit#(8)) ram <- mkRegFileFullLoad("rom.rmh"); // XXX: Make a parameter
    RWire#(Bit#(8)) data_out <- mkRWire;
    TriState#(Bit#(8)) data_tri <- mkTriState(isValid(data_out.wget()), fromMaybe(?, data_out.wget()));

    method Action init_test(MemoryInitT minit);
        for (Integer i=0;i<length(minit);i=i+1) begin
            MemoryInitRunT run = minit[i];
            for (Integer j=0;j<length(run.payload);j=j+1) begin
                ram.upd((run.startaddr + fromInteger(j))[13:0], run.payload[j]);
            end
        end
    endmethod

    // control
    method Action cs(Bit#(1) c);
        cs_in <= c;
    endmethod

    method Action n_oe(Bit#(1) o);
        n_oe_in <= o;
    endmethod

    method Action n_ce(Bit#(1) c);
        n_ce_in <= c;
    endmethod

    // address bus
    method Action addr(Bit#(14) a);
        data_out.wset(ram.sub(a));
    endmethod

    // data bus
    interface data = data_tri.io;
endmodule

endpackage
